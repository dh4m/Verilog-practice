module full_adder (S, A, B, Cout, Cin);

	input A, B, Cin;
	output S, Cout;

// your code

endmodule