module half_adder (S, A, B, C);

	input A, B;
	output S, C;

// your code

endmodule