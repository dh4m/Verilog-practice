`timescale 1ns/100ps

module tb_rca_40b;

// your code

endmodule