module tb_rca_40b;

// your code

endmodule